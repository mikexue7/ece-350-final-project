`timescale 1ns / 1ps
/**
 *
 * READ THIS DESCRIPTION:
 *
 * This is the Wrapper module that will serve as the header file combining your processor,
 * RegFile and Memory elements together.
 *
 * This file will be used to generate the bitstream to upload to the FPGA.
 * We have provided a sibling file, Wrapper_tb.v so that you can test your processor's functionality.
 *
 * We will be using our own separate Wrapper_tb.v to test your code. You are allowed to make changes to the Wrapper files
 * for your own individual testing, but we expect your final processor.v and memory modules to work with the
 * provided Wrapper interface.
 *
 * Refer to Lab 5 documents for detailed instructions on how to interface
 * with the memory elements. Each imem and dmem modules will take 12-bit
 * addresses and will allow for storing of 32-bit values at each address.
 * Each memory module should receive a single clock. At which edges, is
 * purely a design choice (and thereby up to you).
 *
 * You must change line 36 to add the memory file of the test you created using the assembler
 * For example, you would add sample inside of the quotes on line 38 after assembling sample.s
 *
 **/

module Wrapper (clock, reset, up, down, left, right, micData, VGA_R, VGA_G, VGA_B, whichLED, LED_out, hSync, vSync,
	ps2_clk,
  ps2_data,
	reg1, sf,
	chSel, audioOut, audioEn, micClk
	);

	input clock, reset, up, down, left, right, micData;

	inout ps2_clk, ps2_data;


	wire rwe, mwe;
	wire[4:0] rd, rs1, rs2;
	wire[31:0] instAddr, instData,
		rData, regA, regB,
		memAddr, memDataIn, memDataOut;


	output chSel, audioOut, audioEn, micClk;
	output [3:0] VGA_R, VGA_G, VGA_B;
	output [7:0] whichLED;
	output [6:0] LED_out;
	output hSync, vSync;
	output [14:0] reg1;
	output sf;

	wire [5:0] score;
	wire score_flag, isEaten;

	// ADD YOUR MEMORY FILE HERE
	localparam INSTR_FILE = "D:/alternateC/snake_processor/Test Files/Memory Files/addScore";

	// Main Processing Unit
	processor CPU(.clock(clock), .reset(reset),

		// ROM
		.address_imem(instAddr), .q_imem(instData),

		// Regfile
		.ctrl_writeEnable(rwe),     .ctrl_writeReg(rd),
		.ctrl_readRegA(rs1),     .ctrl_readRegB(rs2),
		.data_writeReg(rData), .data_readRegA(regA), .data_readRegB(regB),

		// RAM
		.wren(mwe), .address_dmem(memAddr),
		.data(memDataIn), .q_dmem(memDataOut));

	VGAController Screen(clock, reset, up, left, down, right, score, score_flag, isEaten, hSync, vSync, VGA_R, VGA_G, VGA_B,
			whichLED, LED_out, ps2_clk, ps2_data);

	AudioController A(clock, micData, score_flag, isEaten, chSel, audioOut);

	// Instruction Memory (ROM)
	ROM #(.MEMFILE({INSTR_FILE, ".mem"}))
	InstMem(.clk(clock),
		.addr(instAddr[11:0]),
		.dataOut(instData));

	// Register File
	regfile RegisterFile(.clock(clock),
		.ctrl_writeEnable(rwe), .ctrl_reset(reset),
		.ctrl_writeReg(rd),
		.ctrl_readRegA(rs1), .ctrl_readRegB(rs2),
		.data_writeReg(rData), .data_readRegA(regA), .data_readRegB(regB),
		.score_flag(score_flag), .score(score), .reg1(reg1));

	// Processor Memory (RAM)
	RAM ProcMem(.clk(clock),
		.wEn(mwe),
		.addr(memAddr[11:0]),
		.dataIn(memDataIn),
		.dataOut(memDataOut));

	assign sf = score_flag;
	assign audioEn = 1'b1;

endmodule
